`ifndef BASIC_SYSTEM_SV
    `define BASIC_SYSTEM_SV



`endif 